module EEE_IMGPROC(
	// global clock & reset
	clk,
	reset_n,
	
	// mm slave
	s_chipselect,
	s_read,
	s_write,
	s_readdata,
	s_writedata,
	s_address,

	// stream sink
	sink_data,
	sink_valid,
	sink_ready,
	sink_sop,
	sink_eop,
	
	// streaming source
	source_data,
	source_valid,
	source_ready,
	source_sop,
	source_eop,
	
	// conduit
	mode
	
);


// global clock & reset
input	clk;
input	reset_n;

// mm slave
input							s_chipselect;
input							s_read;
input							s_write;
output	reg	[31:0]	s_readdata;
input	[31:0]				s_writedata;
input	[2:0]					s_address;


// streaming sink
input	[23:0]            	sink_data;
input								sink_valid;
output							sink_ready;
input								sink_sop;
input								sink_eop;

// streaming source
output	[23:0]			  	   source_data;
output								source_valid;
input									source_ready;
output								source_sop;
output								source_eop;

// conduit export
input                         mode;

////////////////////////////////////////////////////////////////////////
//
parameter IMAGE_W = 11'd640;
parameter IMAGE_H = 11'd480;
parameter MESSAGE_BUF_MAX = 256;
parameter MSG_INTERVAL = 6;
parameter BB_COL_DEFAULT = 24'h00ff00;


reg [7:0]   red, green, blue;
wire [7:0]   grey;
wire [7:0]   red_sel, green_sel, blue_sel;

wire [7:0]   red_out, green_out, blue_out;

wire         sop, eop, in_valid, out_ready;
////////////////////////////////////////////////////////////////////////

// Detect red areas
wire tl_detect;
assign tl_detect = red[7] & green[7] & blue[7];

// Find boundary of cursor box

wire [1:0] state;
reg [1:0] next_state;

reg [9:0] x_ctr = 10'b0;
reg [9:0] y_ctr = 10'b0;

assign state = next_state;

// Highlight detected areas
wire [23:0] red_high;
assign grey = green[7:1] + red[7:2] + blue[7:2]; //Grey = green/2 + red/4 + blue/4
assign red_high  =  tl_detect ? {8'hff, 8'hff, 8'hff} : {grey, grey, grey};

// Show bounding box
wire [23:0] new_image;
wire bb_active;
assign bb_active = (x == tl_left) | (x == tl_right) | (y == tl_top) | (y == tl_bottom) | (x == tr_left) | (x == tr_right) | (y == tr_top) | (y == tr_bottom) | (x == bl_left) | (x == bl_right) | (y == bl_top) | (y == bl_bottom) | (x == br_left) | (x == br_right) | (y == br_top) | (y == br_bottom);
assign new_image = bb_active ? bb_col : red_high;

// Switch output pixels depending on mode switch
// Don't modify the start-of-packet word - it's a packet discriptor
// Don't modify data in non-video packets
assign {red_out, green_out, blue_out} = (mode & ~sop & packet_video) ? new_image : {red,green,blue};

//Count valid pixels to tget the image coordinates. Reset and detect packet type on Start of Packet.
reg [10:0] x, y;
reg packet_video;
always@(posedge clk) begin
	if (sop) begin
		x <= 11'h0;
		y <= 11'h0;
		packet_video <= (blue[3:0] == 3'h0);
	end
	else if (in_valid) begin
		if (x == IMAGE_W-1) begin
			x <= 11'h0;
			y <= y + 11'h1;
		end
		else begin
			x <= x + 11'h1;
		end
	end
end

// reg exceeds;

// always begin
// 	if ((x_min == 320) & (x_max == 320) & (y_min ==240) & (y_max == 240)) begin
// 		exceeds = 1;
// 	end
// 	else begin
// 		exceeds = 0;
// 	end
// end
//Find first and last red pixels
reg [10:0] tl_x_min, tl_y_min, tl_x_max, tl_y_max;
reg [10:0] tr_x_min, tr_y_min, tr_x_max, tr_y_max;
reg [10:0] bl_x_min, bl_y_min, bl_x_max, bl_y_max;
reg [10:0] br_x_min, br_y_min, br_x_max, br_y_max;

reg tl_activate, tr_activate, bl_activate, br_activate;

always begin
	if(x >= 320 || y >= 240) begin
		tl_activate = 0;
	end
	else begin
		tl_activate = 1;
	end

	if(x < 320 || y >= 240) begin
		tr_activate = 0;
	end
	else begin
		tr_activate = 1;
	end

	if(x >= 320 || y < 240) begin
		bl_activate = 0;
	end
	else begin
		bl_activate = 1;
	end

	if(x < 320 || y < 240) begin
		br_activate = 0;
	end
	else begin
		br_activate = 1;
	end
end

always@(posedge clk) begin
	if (tl_detect & in_valid & tl_activate) begin	//Update bounds when the pixel is red  & (exceeds == 1'b0)
		if((x < 320) & (x < tl_x_min)) begin
			tl_x_min <= x;
		end
		if((x < 320) & (x > tl_x_max)) begin
			tl_x_max <= x;
		end
		if((y < 240) & (y < tl_y_min)) begin
			tl_y_min <= y;
		end
		if(y < 240) begin
			tl_y_max <= y;
		end
	end

	if (tl_detect & in_valid & tr_activate) begin	//Update bounds when the pixel is red  & (exceeds == 1'b0)
		if((x >= 320) & (x < tr_x_min)) begin
			tr_x_min <= x;
		end
		if((x >= 320) & (x > tr_x_max)) begin
			tr_x_max <= x;
		end
		if((y < 240) & (y < tr_y_min)) begin
			tr_y_min <= y;
		end
		if(y < 240) begin
			tr_y_max <= y;
		end
	end

	if (tl_detect & in_valid & bl_activate) begin	//Update bounds when the pixel is red  & (exceeds == 1'b0)
		if((x < 320) & (x < bl_x_min)) begin
			bl_x_min <= x;
		end
		if((x < 320) & (x > bl_x_max)) begin
			bl_x_max <= x;
		end
		if((y >= 240) & (y < bl_y_min)) begin
			bl_y_min <= y;
		end
		if(y >= 240) begin
			bl_y_max <= y;
		end
	end

	if (tl_detect & in_valid & br_activate) begin	//Update bounds when the pixel is red  & (exceeds == 1'b0)
		if((x >= 320) & (x < br_x_min)) begin
			br_x_min <= x;
		end
		if((x >= 320) & (x > br_x_max)) begin
			br_x_max <= x;
		end
		if((y >= 240) & (y < br_y_min)) begin
			br_y_min <= y;
		end
		if(y >= 240) begin
			br_y_max <= y;
		end
	end

	if (sop & in_valid) begin	//Reset bounds on start of packet
		tl_x_min <= IMAGE_W-11'h1;
		tl_x_max <= 0;
		tl_y_min <= IMAGE_H-11'h1;
		tl_y_max <= 0;

		tr_x_min <= IMAGE_W-11'h1;
		tr_x_max <= 0;
		tr_y_min <= IMAGE_H-11'h1;
		tr_y_max <= 0;

		bl_x_min <= IMAGE_W-11'h1;
		bl_x_max <= 0;
		bl_y_min <= IMAGE_H-11'h1;
		bl_y_max <= 0;

		br_x_min <= IMAGE_W-11'h1;
		br_x_max <= 0;
		br_y_min <= IMAGE_H-11'h1;
		br_y_max <= 0;
	end
end

//Process bounding box at the end of the frame.
reg [1:0] msg_state;
reg [10:0] tl_left, tl_right, tl_top, tl_bottom;
reg [10:0] tr_left, tr_right, tr_top, tr_bottom;
reg [10:0] bl_left, bl_right, bl_top, bl_bottom;
reg [10:0] br_left, br_right, br_top, br_bottom;

reg [7:0] frame_count;
always@(posedge clk) begin
	if (eop & in_valid & packet_video) begin  //Ignore non-video packets
		
		//Latch edges for display overlay on next frame
		tl_left <= tl_x_min;
		tl_right <= tl_x_max;
		tl_top <= tl_y_min;
		tl_bottom <= tl_y_max;

		//Latch edges for display overlay on next frame TR
		tr_left <= tr_x_min;
		tr_right <= tr_x_max;
		tr_top <= tr_y_min;
		tr_bottom <= tr_y_max;

		//Latch edges for display overlay on next frame
		bl_left <= bl_x_min;
		bl_right <= bl_x_max;
		bl_top <= bl_y_min;
		bl_bottom <= bl_y_max;

		//Latch edges for display overlay on next frame TR
		br_left <= br_x_min;
		br_right <= br_x_max;
		br_top <= br_y_min;
		br_bottom <= br_y_max;
		
		//Start message writer FSM once every MSG_INTERVAL frames, if there is room in the FIFO
		frame_count <= frame_count - 1;
		
		if (frame_count == 0 && msg_buf_size < MESSAGE_BUF_MAX - 3) begin
			msg_state <= 2'b01;
			frame_count <= MSG_INTERVAL-1;
		end
	end
	
	//Cycle through message writer states once started
	if (msg_state != 2'b00) msg_state <= msg_state + 2'b01;

end
	

//TODO GENERATE OUTPUT MESSAGES
//Generate output messages for CPU
reg [31:0] msg_buf_in; 
wire [31:0] msg_buf_out;
reg msg_buf_wr;
wire msg_buf_rd, msg_buf_flush;
wire [7:0] msg_buf_size;
wire msg_buf_empty;

`define RED_BOX_MSG_ID "RBB"

always@(*) begin	//Write words to FIFO as state machine advances TODO:ADD NEW BOX HERE
	case(msg_state)
		2'b00: begin
			msg_buf_in = 32'b0;
			msg_buf_wr = 1'b0;
		end
		2'b01: begin
			msg_buf_in = "TL TR BL BR";	//Message ID
			msg_buf_wr = 1'b1;
		end
		2'b10: begin
			msg_buf_in = {tl_x_min, tl_y_min, tr_x_min, tr_y_min, bl_x_min, bl_y_min, br_x_min, br_y_min};	//Top left coordinate
			msg_buf_wr = 1'b1;
		end
		2'b11: begin
			msg_buf_in = {tl_x_max, tl_y_max, tr_x_max, tr_y_max, bl_x_max, bl_y_max, br_x_max, br_y_max}; //Bottom right coordinate
			msg_buf_wr = 1'b1;
		end
	endcase
end



//Output message FIFO
MSG_FIFO	MSG_FIFO_inst (
	.clock (clk),
	.data (msg_buf_in),
	.rdreq (msg_buf_rd),
	.sclr (~reset_n | msg_buf_flush),
	.wrreq (msg_buf_wr),
	.q (msg_buf_out),
	.usedw (msg_buf_size),
	.empty (msg_buf_empty)
);


//Streaming registers to buffer video signal
STREAM_REG #(.DATA_WIDTH(26)) in_reg (
	.clk(clk),
	.rst_n(reset_n),
	.ready_out(sink_ready),
	.valid_out(in_valid),
	.data_out({red,green,blue,sop,eop}),
	.ready_in(out_ready),
	.valid_in(sink_valid),
	.data_in({sink_data,sink_sop,sink_eop})
);

STREAM_REG #(.DATA_WIDTH(26)) out_reg (
	.clk(clk),
	.rst_n(reset_n),
	.ready_out(out_ready),
	.valid_out(source_valid),
	.data_out({source_data,source_sop,source_eop}),
	.ready_in(source_ready),
	.valid_in(in_valid),
	.data_in({red_out, green_out, blue_out, sop, eop})
);


/////////////////////////////////
/// Memory-mapped port		 /////
/////////////////////////////////

// Addresses
`define REG_STATUS    			0
`define READ_MSG    				1
`define READ_ID    				2
`define REG_BBCOL					3

//Status register bits
// 31:16 - unimplemented
// 15:8 - number of words in message buffer (read only)
// 7:5 - unused
// 4 - flush message buffer (write only - read as 0)
// 3:0 - unused


// Process write

reg  [7:0]   reg_status;
reg	[23:0]	bb_col;

always @ (posedge clk)
begin
	if (~reset_n)
	begin
		reg_status <= 8'b0;
		bb_col <= BB_COL_DEFAULT;
	end
	else begin
		if(s_chipselect & s_write) begin
		   if      (s_address == `REG_STATUS)	reg_status <= s_writedata[7:0];
		   if      (s_address == `REG_BBCOL)	bb_col <= s_writedata[23:0];
		end
	end
end


//Flush the message buffer if 1 is written to status register bit 4
assign msg_buf_flush = (s_chipselect & s_write & (s_address == `REG_STATUS) & s_writedata[4]);


// Process reads
reg read_d; //Store the read signal for correct updating of the message buffer

// Copy the requested word to the output port when there is a read.
always @ (posedge clk)
begin
   if (~reset_n) begin
	   s_readdata <= {32'b0};
		read_d <= 1'b0;
	end
	
	else if (s_chipselect & s_read) begin
		if   (s_address == `REG_STATUS) s_readdata <= {16'b0,msg_buf_size,reg_status};
		if   (s_address == `READ_MSG) s_readdata <= {msg_buf_out};
		if   (s_address == `READ_ID) s_readdata <= 32'h1234EEE2;
		if   (s_address == `REG_BBCOL) s_readdata <= {8'h0, bb_col};
	end
	
	read_d <= s_read;
end

//Fetch next word from message buffer after read from READ_MSG
assign msg_buf_rd = s_chipselect & s_read & ~read_d & ~msg_buf_empty & (s_address == `READ_MSG);
						


endmodule

